* C:\Pooja hacakathon\LDO.cir

*** Spice lib***

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

******* Transistor Connection*****
xM4   net_d    Vb4     net3     GND  sky130_fd_pr__nfet_01v8
xM2   net1     net_d   VDD      VDD  sky130_fd_pr__pfet_01v8
xM1   net3     net_R2  net_diff GND  sky130_fd_pr__nfet_01v8
xM44  Vgpass   Vb4     net4     GND  sky130_fd_pr__nfet_01v8
xM11  net4     VREF    net_diff GND  sky130_fd_pr__nfet_01v8
xM3   net_d    Vb3     net1     VDD  sky130_fd_pr__pfet_01v8
xM33  Vgpass   Vb3     net2     VDD  sky130_fd_pr__pfet_01v8
xM55  net_diff VDD     GND      GND  sky130_fd_pr__nfet_01v8
xM5   VDD      VDD     GND      GND  sky130_fd_pr__nfet_01v8
xMP1  Vout     Vgpass  VDD      VDD  sky130_fd_pr__pfet_01v8
xM02  GND      GND     net_d1   VDD  sky130_fd_pr__pfet_01v8
xM0   net_R2   net_R2  Vout     VDD  sky130_fd_pr__pfet_01v8
xM01  net_d1   net_d1  net_R2   VDD  sky130_fd_pr__pfet_01v8
xM22  net2     net_d   VDD      VDD  sky130_fd_pr__pfet_01v8
C2    Vout     GND     1p


***** Power Potential*******

Vdd vdd 0 3.3
Vb3 vb3 0 0
Vb4 vb4 0 3.3
VREF VREF 0 1.2

**** Analysis*****

*.tran 5e-09 20e-09 0e-09

.dc vdd 2e-00 3.3e-00 0.1e-00

* Control Statements

.control
run

**** Output Plot****

plot V(vdd) V(Vout)
plot V(Vout) vs V(Vdd)

.endc
.end
